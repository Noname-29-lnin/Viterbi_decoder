module tb_Testcase2();

endmodule
