module viterbi_deocode(
   input logic          i_clk,
   input logic          i_rst_n,

   input logic [1:0]    i_input_data,

   output logic         o_output_data
);
// Wire
wire w_done;
wire [1:0] w_input_data;
wire [1:0] w_BM_0, w_BM_1, w_BM_2, w_BM_3;
wire [1:0] w_iPM_0, w_iPM_1, w_iPM_2, w_iPM_3;
wire [1:0] w_oPM_0, w_oPM_1, w_oPM_2, w_oPM_3;

d_ff DFF_BMU(
    .i_clk      (i_clk),
    .i_rst_n    (i_rst_n),
    .i_en       (w_done),
    .i_data     (i_input_data),
    .o_data     (w_input_data)
);
branch_metric_unit  BMU(
    // input logic         i_clk,
    // input logic         i_rst_n,
    // input logic         i_en,
    .i_data             (w_input_data),
    .o_branch_metric_0  (w_BM_0),
    .o_branch_metric_1  (w_BM_1),
    .o_branch_metric_2  (w_BM_2),
    .o_branch_metric_3  (w_BM_3)
);
Add_compare_select_unit ACSU(
    // input logic     i_clk,
    // input logic     i_rst_n,
    // input logic     i_en,

    .i_branch_metric_0      (w_BM_0),
    .i_branch_metric_1      (w_BM_1),
    .i_branch_metric_2      (w_BM_2),
    .i_branch_metric_3      (w_BM_3),

    .i_path_metric_0        (w_iPM_0),
    .i_path_metric_1        (w_iPM_1),
    .i_path_metric_2        (w_iPM_2),
    .i_path_metric_3        (w_iPM_3),

    .o_path_metric_0        (w_oPM_0),
    .o_path_metric_1        (w_oPM_1),
    .o_path_metric_2        (w_oPM_2),
    .o_path_metric_3        (w_oPM_3)

    // output logic       o_done
);
path_metric_unit PMU(
    .i_clk                  (i_clk),
    .i_rst_n                (i_rst_n),
    .i_en                   (w_done),

    .i_path_metric_0        (w_oPM_0),
    .i_path_metric_1        (w_oPM_1),
    .i_path_metric_2        (w_oPM_2),
    .i_path_metric_3        (w_oPM_3),

    .o_path_metric_0        (w_iPM_0),
    .o_path_metric_1        (w_iPM_1),
    .o_path_metric_2        (w_iPM_2),
    .o_path_metric_3        (w_iPM_3)
);
survivor_path_memory SPMU(
    .i_clk              (i_clk),
    .i_rst_n            (i_rst_n),
    .i_path_metric_0    (w_oPM_0),
    .i_path_metric_1    (w_oPM_1),
    .i_path_metric_2    (w_oPM_2), 
    .i_path_metric_3    (w_oPM_3),
    
    .o_decision_bit     (o_output_data),
    .o_done             (w_done)
);

endmodule