module Add_unit(
    input logic [1:0]       i_BM    ,
    input logic [1:0]       i_PM    ,
    output logic [1:0]      o_PM    
);

// | A  | B  | S  |
// | 00 | 00 | 00 |
// | 00 | 01 | 01 |
// | 00 | 10 | 10 |
// | 00 | 11 | 11 |
// | 01 | 00 | 01 |
// | 01 | 01 | 10 |
// | 01 | 10 | 11 |
// | 01 | 11 | 11 |
// | 10 | 00 | 10 |
// | 10 | 01 | 11 |
// | 10 | 10 | 11 |
// | 10 | 11 | 11 |
// | 11 | 00 | 11 |
// | 11 | 01 | 11 |
// | 11 | 10 | 11 |
// | 11 | 11 | 11 |

assign o_PM[0] = (!i_PM[0]&i_BM[0]) | (i_PM[0]&!i_BM[0]) | 
                 (i_PM[0]&i_BM[1]) | (i_PM[1]&i_BM[0])   | 
                 (i_PM[1]&i_BM[1]);
assign o_PM[1] = (i_PM[1] | i_BM[1]) | (i_PM[0] & i_BM[0]);

endmodule
